
//------------------------------------------------------------------------------
// apb transfer enums, parameters, and events
typedef enum { APB_READ = 0, APB_WRITE = 1 } apb_direction_enum;
